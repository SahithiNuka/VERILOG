module mux_10x1_tb();
	reg [9:0]i;
	reg [3:0]s;
	wire y;
	
	mux_10x1 m1(i,s,y);
	
	initial
		begin
			i = 10'b1010101011;
			s = 4'd0;
			#10;
			
			i = 10'b1010101011;
			s = 4'd1;
			#10;
			
			i = 10'b1010101011;
			s = 4'd2;
			#10;
			
			i = 10'b1010101011;
			s = 4'd3;
			#10;
			
			i = 10'b1010101011;
			s = 4'd4;
			#10;
			
			i = 10'b1010101011;
			s = 4'd5;
			#10;
			
			i = 10'b1010101011;
			s = 4'd6;
			#10;
			
			i = 10'b1010101011;
			s = 4'd7;
			#10;
			
			i = 10'b1010101011;
			s = 4'd8;
			#10;
			
			i = 10'b1010101011;
			s = 4'd9;
			#10;
			
			i = 10'b1010101011;
			s = 4'd10;
			#10;
			
			i = 10'b1010101011;
			s = 4'd11;
			#10;
			
			i = 10'b1010101011;
			s = 4'd12;
			#10;
			
			i = 10'b1010101011;
			s = 4'd13;
			#10;
			
			i = 10'b1010101011;
			s = 4'd14;
			#10;
			
			i = 10'b1010101011;
			s = 4'd15;
			#10;
			$finish;
		end
		
		initial
			$monitor("i=%b,s=%b,y=%b",i,s,y);
endmodule