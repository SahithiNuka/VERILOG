module seq_detector_10010_mealy_2bit_overlapping_tb();
	reg clk;
	reg reset;
	reg din;
	wire dout;
	
  	seq_detector_10010_mealy_2bit_overlapping uut (clk,reset,din,dout);
	
	initial
		begin
			clk=1'b1;
			forever #5 clk = ~clk;
		end
	
	// Task to apply one bit input in sync with clock 
	task apply_bit(input value);
		begin
			@(negedge clk);
			din = value;
			@(posedge clk); // wait for clock positive edge to latch
		end
	endtask
	
	initial begin
		reset = 1;
		din = 0;
		#15;
		reset = 0;
		
		// Apply input bits with interval of one clock cycle
		// Sequence: 10010 (should detect)
		apply_bit(1);
		apply_bit(0);
		apply_bit(0);
		apply_bit(1);
		apply_bit(0);
		
		// Random bits no detection
		apply_bit(1);
		apply_bit(0);
		apply_bit(0);
		apply_bit(1);
		apply_bit(1);
		
		// Some random bits to show 2-bit overlapping behavior
		apply_bit(1);
		apply_bit(0);
		apply_bit(0);
		apply_bit(1);
		apply_bit(0);
		
		apply_bit(0);
		apply_bit(1);
		apply_bit(0);
		
		#20;
		$finish;
	end

	initial begin
		$monitor("t=%t, reset=%b, din=%b, dout=%b",$time,reset,din,dout);
	end
  
	initial
		begin
			$dumpfile("dump.vcd");
			$dumpvars;
		end

endmodule